
module address_change (
